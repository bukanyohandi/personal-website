`timescale 1ns/1ps
`include "ALU.v"

module alu_test;

reg[31:0] instruction, regA, regB;

wire[31:0] result;
wire[2:0] flags;

alu test_ALU(instruction, regA, regB, result, flags);

initial
    begin

    $display("instruction:op:func:  regA  :  regB  :   rs   :   rt   : result :z:n:o");
    $monitor("   %h:%h: %h :%h:%h:%h:%h:%h:%h:%h:%h",
    instruction, test_ALU.opcode, test_ALU.func, regA, regB, test_ALU.rs, test_ALU.rt, result, flags[2], flags[1], flags[0]);

    // [1] add $t0 regA regB, expect: overflow flag
    #10 instruction <= 32'b0000_0000_0000_0001_0100_0000_0010_0000;
    regA <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;
    regB <= 32'b0100_0000_0000_0000_0000_0000_0000_0000;

    // [2] addi $t1 regA 13 
    #10 instruction <= 32'b0010_0000_0000_1001_0000_0000_0000_1101;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;

    // [3] addu $t2 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0101_0000_0010_0001;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1001;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0100;

    // [4] addiu $t3 regA 13 
    #10 instruction <= 32'b0010_0100_0000_1011_0000_0000_0000_1101;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0011;

    // [5] sub $t0 regA regB, expect: overflow flag
    #10 instruction <= 32'b0000_0000_0000_0001_0100_0000_0010_0010;
    regA <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0001;

    // [6] subu $t1 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0100_1000_0010_0011;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;

    // [7] and $t0 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0100_0000_0010_0100;
    regA <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
    regB <= 32'b0000_0000_0000_0000_0110_0111_1001_1000;

    // [8] andi $t1 regA 13 
    #10 instruction <= 32'b0011_0000_0000_1001_0000_0000_0000_1101;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;

    // [9] nor $t2 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0101_0000_0010_0111;
    regA <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
    regB <= 32'b0110_1001_0110_1001_0110_1001_0110_1001;

    // [10] or $t3 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0101_1000_0010_0101;
    regA <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
    regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;

    // [11] ori $t4 regA 13 
    #10 instruction <= 32'b0011_0100_0000_1100_0000_0000_0000_1101;
    regA <= 32'b0000_0000_0000_0000_0000_0001_1000_0010;

    // [12] xor $t5 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0110_1000_0010_0110;
    regA <= 32'b1000_0111_0110_0101_0100_0011_0010_0001;
    regB <= 32'b0001_0010_0011_0100_0101_0110_0111_1000;

    // [13] xori $t6 regA 13 
    #10 instruction <= 32'b0011_1000_0000_1110_0000_0000_0000_1101;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0101_0100;

    // [14] beq regA regB 13 
    #10 instruction <= 32'b0001_0000_0000_0001_1111_1111_1111_1111;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;

    // [15] bne regA regB 13, expect: zero flag 
    #10 instruction <= 32'b0001_0100_0000_0001_1111_1111_1111_1111;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0110;

    // [16] slt $t0 regA regB 
    #10 instruction <= 32'b0000_0000_0000_0001_0100_0000_0010_1010;
    regA <= 32'b0000_0000_0000_0000_1111_1110_1100_1000;
    regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;

    // [17] slti $t1 regA 13, expect: negative flag
    #10 instruction <= 32'b0010_1000_0000_1001_0000_0000_0000_1101;
    regA <= 32'b1000_0000_0000_0000_0000_0000_0000_1000;

    // [18] sltiu $t2 regA 13 
    #10 instruction <= 32'b0010_1100_0000_1010_0000_0000_0000_1101;
    regA <= 32'b1000_0000_0000_0000_0000_0000_0000_1000;

    // [19] sltu $t3 regA regB, expect: negative flag
    #10 instruction <= 32'b0000_0000_0000_0001_0101_1000_0010_1011;
    regA <= 32'b0000_0000_0000_0000_1111_1110_1100_1000;
    regB <= 32'b1000_0000_0000_0000_0000_0000_0000_0000;

    // [20] lw $t1 1(regB) 
    #10 instruction <= 32'b1000_1100_0010_1001_0000_0000_0000_0001;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_1110;

    // [21] sw $t2 1(regA) 
    #10 instruction <= 32'b1010_1100_0000_1010_0000_0000_0000_0001;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1110;

    // [22] sll $t0 regA 13 
    #10 instruction <= 32'b0000_0000_0000_0000_0100_0011_0100_0000;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;

    // [23] sllv $t1 regA regB 
    #10 instruction <= 32'b0000_0000_0010_0000_0100_1000_0000_0100;
    regA <= 32'b0000_0000_0000_0000_0000_0000_0000_1111;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_1101;

    // [24] srl $t2 regA 13 
    #10 instruction <= 32'b0000_0000_0000_0000_0101_0011_0100_0010;
    regA <= 32'b1000_1100_1110_0000_0000_0000_0000_0000;

    // [25] srlv $t3 regA regB 
    #10 instruction <= 32'b0000_0000_0010_0000_0101_1000_0000_0110;
    regA <= 32'b0010_0110_0001_0101_1000_0000_0000_0000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_0101;

    // [26] sra $t4 regA 13 
    #10 instruction <= 32'b0000_0000_0000_0000_0110_0011_0100_0011;
    regA <= 32'b1110_1010_0110_0001_1000_0000_0000_0000;

    // [27] srav $t5 regA regB 
    #10 instruction <= 32'b0000_0000_0010_0000_0110_1000_0000_0111;
    regA <= 32'b1110_1010_0110_0001_1000_0000_0000_0000;
    regB <= 32'b0000_0000_0000_0000_0000_0000_0000_1101;

    #10 $finish;
    end
endmodule